// unnamed.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module unnamed (
		input  wire        address,    //  avalon_irda_slave.address
		input  wire        chipselect, //                   .chipselect
		input  wire [3:0]  byteenable, //                   .byteenable
		input  wire        read,       //                   .read
		input  wire        write,      //                   .write
		input  wire [31:0] writedata,  //                   .writedata
		output wire [31:0] readdata,   //                   .readdata
		input  wire        clk,        //                clk.clk
		output wire        IRDA_TXD,   // external_interface.TXD
		input  wire        IRDA_RXD,   //                   .RXD
		output wire        irq,        //          interrupt.irq
		input  wire        reset       //              reset.reset
	);

	unnamed_irda_0 irda_0 (
		.clk        (clk),        //                clk.clk
		.reset      (reset),      //              reset.reset
		.address    (address),    //  avalon_irda_slave.address
		.chipselect (chipselect), //                   .chipselect
		.byteenable (byteenable), //                   .byteenable
		.read       (read),       //                   .read
		.write      (write),      //                   .write
		.writedata  (writedata),  //                   .writedata
		.readdata   (readdata),   //                   .readdata
		.irq        (irq),        //          interrupt.irq
		.IRDA_TXD   (IRDA_TXD),   // external_interface.export
		.IRDA_RXD   (IRDA_RXD)    //                   .export
	);

endmodule
