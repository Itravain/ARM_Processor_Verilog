module tester(
	input wire [31:0] entrada_um, entrada_dois,
	output wire [31:0] saida_um, saida_dois
);
	
	assign saida_um = entrada_um;
	assign saida_dois = entrada_dois;

endmodule 